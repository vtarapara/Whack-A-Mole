`timescale 1 ns / 100 ps

module regfile_tb();
    
endmodule
